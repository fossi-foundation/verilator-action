module B;
    wire [1:0] b;

    assign b = 1'b1;
endmodule