module A;
    wire [1:0] a;

    assign a = 1'b1;
endmodule